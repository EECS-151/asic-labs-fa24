module shift_register_behavioral (
    input in,
    input clk,
    output [3:0] out
);
    reg [3:0] shift_reg;

    always @(posedge clk) begin
        // TODO
    end

    ____ out = ____; // TODO
endmodule
